`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/07/2023 02:20:43 PM
// Design Name: 
// Module Name: Hazard_Detection_Unit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Hazard_Detection_Unit(
    input [4:0] rs1,
    input [4:0] rs2,
    input de_ex_memRead,
    input [4:0] de_ex_regRd,
    output logic de_write,
    output logic pcWrite,
    output logic controlMux,
    output logic loadUse,
    output logic branchValid
    );
    
    
    
    
endmodule
